module b;
endmodule
