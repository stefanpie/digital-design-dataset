module a;
b b_inst ();
c c_inst ();
endmodule
