module d;
endmodule
