module b;
endmodule

module c;
d d_inst ();
endmodule
