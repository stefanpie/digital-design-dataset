module c;
endmodule
