module a;
b b_inst ();
c c_inst ();
endmodule

module a_prime;
b b_inst ();
c c_inst ();
endmodule

module b;
endmodule

module c;
endmodule

